module gas_csr (
    input wire i_sig_csrr,
    input wire [1:0] i_csrr,
    input wire [11:0] i_csr_addr,

    output wire [63:0] o_csr_data
);
    
endmodule