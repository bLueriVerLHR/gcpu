module gf_if #(
    ADDR_LEN  = 64,
    INST_LEN  = 32,
    INST_BLEN = 4
) (
    input pc
);
endmodule